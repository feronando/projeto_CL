library verilog;
use verilog.vl_types.all;
entity projeto_CL_vlg_vec_tst is
end projeto_CL_vlg_vec_tst;
